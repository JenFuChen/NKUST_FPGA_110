library verilog;
use verilog.vl_types.all;
entity HW_vlg_vec_tst is
end HW_vlg_vec_tst;
