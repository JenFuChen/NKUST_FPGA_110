module HW2(CLK,en,count);
input CLK,en ; 
output [3:0] count; 
reg [3:0] count; 
always@(posedge CLK)
begin 
if(!en) 
count<=8'h0; //nonblocking 
else 
if(count==8'h9)
	count=0;
else
	count<=count+ 1;
end 
endmodule
