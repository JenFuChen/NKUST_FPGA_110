module hw();
intput  







endmodule
