library verilog;
use verilog.vl_types.all;
entity hw3_vlg_vec_tst is
end hw3_vlg_vec_tst;
